
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity t_flipflop is 
port( 
t,clk ,clr :in std_logic ;
q:out std_logic );
end t_flipflop;

architecture tff of t_flipflop is
signal s:std_logic:='0';
begin 
process (t,clk,clr)
begin
if clr='0' then s<= '0';

elsif rising_edge(clk)then 

if t<='0' then s<=s;
else s<= not (s);

end if;
end if;
end process;
q<= s;
end tff;